// Include all the testbench files here. The order of files is the order in which they compile. 
//`include "./../uvc/fifo_driver.sv"
// include fifo_agent, fifo_env and fifo_test files in the order it is mentioned.  

`include "./../test/msg_test.sv"


